// my_macros.vh - placeholder macros file

`define MY_MACRO 1
